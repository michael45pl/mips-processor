library IEEE;
use IEEE.std_logic_1164.all;

entity control is
  port( func : in std_logic_vector(5 downto 0);
	op   : in std_logic_vector(5 downto 0);
	ALUControl 	: out std_logic_vector(5 downto 0);
	ALUSrc    	: out std_logic;
	ALU_shift    	: out std_logic;
	MemToReg   	: out std_logic;
	RegDst     	: out std_logic;
	s_DMemWr   	: out std_logic;
	s_RegWr    	: out std_logic;
	jump	   	: out std_logic;
	branch		: out std_logic;
	upper		: out std_logic;
	jr		: out std_logic;
	jal		: out std_logic;
	extend		: out std_logic;
	bne		: out std_logic);
end control;

architecture structure of control is

begin

  p_CASE : process (func, op)

  begin

	case op is
      	when "000000" =>
      		case func is
      		when "100000" => --add
      			ALUControl <= "000110"; -- x6 is add
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when "100001" => --addu
      			ALUControl <= "000110"; -- x6 is add
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when "100100" => --and
      			ALUControl <= "000000"; -- x0 is and
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when "100101" => --or
      			ALUControl <= "000001"; -- x1 is or
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when "100110" => --xor
      			ALUControl <= "000010"; -- x2 is xor
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when "100111" => --nor
      			ALUControl <= "000100"; -- x4 is or
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "101010" => --slt
      			ALUControl <= "000101"; -- x5 is slt
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "101011" => --sltu
      			ALUControl <= "000101"; -- x5 is slt
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000000" => --sll
      			ALUControl <= "000010"; -- x0 is sll
      			ALUSrc     <= '1'; -- uses shamt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '0'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000010" => --srl
      			ALUControl <= "000000"; -- x1 is srl
      			ALUSrc     <= '1'; -- uses shamt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000011" => --sra
      			ALUControl <= "000001"; -- x3 is sra
      			ALUSrc     <= '1'; -- uses shamt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000100" => --sllv
      			ALUControl <= "000010"; -- x0 is sll
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000110" => --srlv
      			ALUControl <= "000000"; -- x2 is srl
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "000111" => --srav
      			ALUControl <= "000001"; -- x3 is sra
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '1'; -- uses shifter so 1
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "100010" => --sub
      			ALUControl <= "000111"; -- x7 is sub
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
          when "100011" => --subu
      			ALUControl <= "000111"; -- x7 is sub
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '1'; -- writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '0'; -- zero extend
			bne	   <= '0'; -- not bne
	when "001000" => --jr
      			ALUControl <= "000000"; -- ?
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '1'; -- writes to rd
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '0'; -- not writing to reg
			jump  	   <= '0'; -- jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '1'; -- is jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		when others =>
      			ALUControl <= "000000"; -- x0 is and
      			ALUSrc     <= '0'; -- uses rt
			ALU_shift  <= '0'; -- uses ALU so 0
      			MemToReg   <= '0'; -- doesn't use mem
      			RegDst     <= '0'; -- writes to rt
      			s_DMemWr   <= '0'; -- not writing to mem
      			s_RegWr    <= '0'; -- not writing to reg
			jump	   <= '0'; -- not jump
			branch	   <= '0'; -- not branch
			upper	   <= '0'; -- not upper
			jr	   <= '0'; -- not jr
			jal	   <= '0'; -- not jal
			extend	   <= '1'; -- sign extend
			bne	   <= '0'; -- not bne
      		end case;
      	when "001000" => --addi
      		ALUControl <= "000110"; -- x6 is add
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
      	when "001001" => --addiu
      		ALUControl <= "000110"; -- x6 is add
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
      	when "001100" => --andi
      		ALUControl <= "000000"; -- x0 is and
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '1'; -- writes to rd
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '0'; -- zero extend
		bne	   <= '0'; -- not bne
      	when "001111" => --lui
      		ALUControl <= "000110"; -- ?
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- ?
      		MemToReg   <= '0'; -- writes from ALU
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '1'; -- is upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
      	when "100011" => --lw
      		ALUControl <= "000110"; -- x6 is add
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '1'; -- writes from mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
      	when "001110" => --xori
      		ALUControl <= "000010"; -- x2 is xor
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '0'; -- zero extend
		bne	   <= '0'; -- not bne
      	when "001101" => --ori
      		ALUControl <= "000001"; -- x1 is or
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '0'; -- zero extend
		bne	   <= '0'; -- not bne
        when "001010" => --slti
      		ALUControl <= "000101"; -- x5 is slt
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
        when "001011" => --sltiu
      		ALUControl <= "000101"; -- x5 is slt
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
        when "101011" => --sw
      		ALUControl <= "000110"; -- x6 is add
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't write from mem
      		RegDst     <= '1'; -- writes to rd
      		s_DMemWr   <= '1'; -- writing to mem
      		s_RegWr    <= '0'; -- not writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
	when "000101" => --bne
      		ALUControl <= "000111"; -- x7 is sub
      		ALUSrc     <= '0'; -- uses rt
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '1'; -- writes to rd
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '0'; -- writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '1'; -- branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- writes to pc like jal ---changed from 1
		extend	   <= '1'; -- sign extend
		bne	   <= '1'; -- is bne
	when "000100" => --beq
      		ALUControl <= "000111"; -- x7 is sub
      		ALUSrc     <= '0'; -- uses rt
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '1'; -- writes to rd
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '0'; -- not writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '1'; -- branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
	when "000010" => --j
      		ALUControl <= "000000"; -- ?
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '1'; -- writes to rd
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '0'; -- not writing to reg
		jump  	   <= '1'; -- jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '0'; -- zero extend
		bne	   <= '0'; -- not bne
	when "000011" => --jal
      		ALUControl <= "000000"; -- ?
      		ALUSrc     <= '1'; -- uses imm
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- doesn't writes to rd
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '1'; -- writing to reg
		jump  	   <= '1'; -- jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '1'; -- is jal
		extend	   <= '0'; -- zero extend
		bne	   <= '0'; -- not bne
      	when others =>
      		ALUControl <= "000000"; -- x0 is and
      		ALUSrc     <= '0'; -- uses rt
		ALU_shift  <= '0'; -- uses ALU so 0
      		MemToReg   <= '0'; -- doesn't use mem
      		RegDst     <= '0'; -- writes to rt
      		s_DMemWr   <= '0'; -- not writing to mem
      		s_RegWr    <= '0'; -- not writing to reg
		jump  	   <= '0'; -- not jump
		branch	   <= '0'; -- not branch
		upper	   <= '0'; -- not upper
		jr	   <= '0'; -- not jr
		jal	   <= '0'; -- not jal
		extend	   <= '1'; -- sign extend
		bne	   <= '0'; -- not bne
    	end case;

  end process;

end structure;
