library IEEE;
use IEEE.std_logic_1164.all;

package regarr is
	type reg_arr is array(0 to 31) of std_logic;
end package regarr;